library ieee;
use ieee.std_logic_1164.all;

entity top is
end top;

architecture behav of top is

begin


end behav;

