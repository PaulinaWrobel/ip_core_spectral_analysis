library ieee;
use ieee.std_logic_1164.all;

entity spectral_analysis is

end entity spectral_analysis;

architecture Behavioral of spectral_analysis is

begin


end architecture Behavioral;

