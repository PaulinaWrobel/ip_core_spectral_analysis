library ieee;
use ieee.std_logic_1164.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

entity top is
end top;

architecture behav of top is

begin


end behav;

